// Actel Corporation Proprietary and Confidential
//  Copyright 2008 Actel Corporation.  All rights reserved.
// ANY USE OR REDISTRIBUTION IN PART OR IN WHOLE MUST BE HANDLED IN
// ACCORDANCE WITH THE ACTEL LICENSE AGREEMENT AND MUST BE APPROVED
// IN ADVANCE IN WRITING.
//  Revision Information:
// Jun09    Revision 4.1
// Aug10    Revision 4.2
// SVN Revision Information:
// SVN $Revision: 8508 $
// SVN $Date: 2009-06-15 16:49:49 -0700 (Mon, 15 Jun 2009) $
`timescale 1ns/1ns
module
COREUART_C0_COREUART_C0_0_COREUART
(
RESET_N
,
CLK
,
WEN
,
OEN
,
CSN
,
DATA_IN
,
RX
,
BAUD_VAL
,
BIT8
,
PARITY_EN
,
ODD_N_EVEN
,
PARITY_ERR
,
OVERFLOW
,
TXRDY
,
RXRDY
,
DATA_OUT
,
TX
,
FRAMING_ERR
,
BAUD_VAL_FRACTION
)
;
parameter
TX_FIFO
=
0
;
parameter
RX_FIFO
=
0
;
parameter
RX_LEGACY_MODE
=
0
;
parameter
FAMILY
=
15
;
parameter
BAUD_VAL_FRCTN_EN
=
0
;
parameter
SYNC_RESET
=
(
FAMILY
==
25
)
?
1
:
0
;
input
RESET_N
;
input
CLK
;
input
WEN
;
input
OEN
;
input
CSN
;
input
[
7
:
0
]
DATA_IN
;
input
RX
;
input
[
12
:
0
]
BAUD_VAL
;
input
BIT8
;
input
PARITY_EN
;
input
ODD_N_EVEN
;
input
[
2
:
0
]
BAUD_VAL_FRACTION
;
output
PARITY_ERR
;
output
OVERFLOW
;
output
TXRDY
;
output
RXRDY
;
output
[
7
:
0
]
DATA_OUT
;
output
TX
;
output
FRAMING_ERR
;
`define CUARTOII  \
2 \
'b \
00
`define CUARTIII  \
2 \
'b \
01
`define CUARTlII  \
2 \
'b \
10
`define CUARTOlI  \
2 \
'b \
11
wire
PARITY_ERR
;
wire
FRAMING_ERR
;
wire
OVERFLOW
;
wire
CUARTIlI
;
wire
TXRDY
;
reg
RXRDY
;
wire
CUARTllI
;
wire
CUARTO0I
;
wire
CUARTI0I
;
reg
[
7
:
0
]
DATA_OUT
;
wire
TX
;
wire
CUARTll
;
wire
CUARTIl
;
wire
CUARTl0I
;
reg
[
7
:
0
]
CUARTO1I
;
wire
[
7
:
0
]
CUARTI1I
;
wire
[
7
:
0
]
CUARTl1I
;
wire
CUARTOOl
;
reg
[
7
:
0
]
CUARTIOl
;
wire
[
7
:
0
]
CUARTlOl
;
wire
[
7
:
0
]
CUARTOIl
;
wire
CUARTIIl
;
wire
CUARTlIl
;
reg
CUARTOll
;
reg
CUARTIll
;
wire
CUARTlll
;
wire
CUARTO0l
;
wire
CUARTI0l
;
wire
CUARTl0l
;
wire
CUARTO1l
;
wire
CUARTI1l
;
reg
CUARTl1l
;
reg
CUARTOO0
;
wire
CUARTIO0
;
reg
CUARTlO0
;
reg
CUARTOI0
;
reg
CUARTII0
;
reg
CUARTlI0
;
reg
CUARTOl0
;
reg
CUARTIl0
;
reg
[
1
:
0
]
CUARTll0
;
reg
[
1
:
0
]
CUARTO00
;
wire
CUARTI00
;
wire
CUARTl00
;
reg
CUARTO10
;
wire
CUARTI10
;
wire
CUARTI1
;
wire
CUARTl1
;
assign
CUARTI1
=
(
SYNC_RESET
==
1
)
?
1
'b
1
:
RESET_N
;
assign
CUARTl1
=
(
SYNC_RESET
==
1
)
?
RESET_N
:
1
'b
1
;
always
@
(
posedge
CLK
or
negedge
CUARTI1
)
begin
:
CUARTl10
if
(
(
!
CUARTI1
)
||
(
!
CUARTl1
)
)
begin
CUARTO1I
<=
{
8
{
1
'b
0
}
}
;
CUARTIll
<=
1
'b
1
;
end
else
begin
CUARTIll
<=
1
'b
1
;
if
(
CSN
==
1
'b
0
&
WEN
==
1
'b
0
)
begin
CUARTO1I
<=
DATA_IN
;
CUARTIll
<=
1
'b
0
;
end
end
end
assign
CUARTl0I
=
WEN
==
1
'b
0
&
CSN
==
1
'b
0
?
1
'b
1
:
1
'b
0
;
always
@
(
CUARTlOl
or
CUARTIOl
or
PARITY_ERR
)
begin
if
(
RX_FIFO
==
1
'b
0
)
begin
DATA_OUT
=
CUARTlOl
;
end
else
begin
if
(
PARITY_ERR
==
1
'b
1
)
begin
DATA_OUT
=
CUARTlOl
;
end
else
begin
DATA_OUT
=
CUARTIOl
;
end
end
end
assign
CUARTOOl
=
(
RX_FIFO
==
1
'b
0
)
?
(
(
CSN
==
1
'b
0
&
OEN
==
1
'b
0
)
?
1
'b
1
:
1
'b
0
)
:
!
CUARTI0l
;
assign
CUARTl0l
=
(
RX_FIFO
==
1
'b
0
)
?
(
(
CSN
==
1
'b
0
&
OEN
==
1
'b
0
)
?
1
'b
1
:
1
'b
0
)
:
CUARTOO0
;
assign
CUARTO1l
=
(
RX_FIFO
==
1
'b
0
)
?
(
(
CSN
==
1
'b
0
&
OEN
==
1
'b
0
)
?
1
'b
1
:
1
'b
0
)
:
(
(
CSN
==
1
'b
0
&
OEN
==
1
'b
0
)
?
1
'b
1
:
CUARTOI0
)
;
assign
CUARTI10
=
(
CSN
==
1
'b
0
&
OEN
==
1
'b
0
)
?
1
'b
1
:
1
'b
0
;
assign
CUARTOIl
=
(
PARITY_ERR
==
1
'b
0
)
?
CUARTlOl
:
8
'b
0
;
generate
if
(
RX_LEGACY_MODE
==
1
'b
1
)
begin
always
@
(
CUARTllI
or
CUARTOl0
)
begin
if
(
RX_FIFO
==
1
'b
0
)
begin
RXRDY
=
CUARTllI
;
end
else
begin
RXRDY
=
!
CUARTOl0
;
end
end
end
else
begin
always
@
(
posedge
CLK
or
negedge
CUARTI1
)
begin
if
(
(
!
CUARTI1
)
||
(
!
CUARTl1
)
)
begin
RXRDY
<=
1
'b
0
;
end
else
begin
if
(
RX_FIFO
==
1
'b
0
)
begin
if
(
CUARTI00
==
1
'b
1
||
CUARTllI
==
1
'b
0
)
begin
RXRDY
<=
CUARTllI
;
end
end
else
begin
if
(
CUARTI00
==
1
'b
1
||
(
CUARTOl0
==
1
'b
1
)
||
(
(
CUARTOl0
==
1
'b
0
)
&&
(
CUARTl00
==
1
'b
1
||
RX_FIFO
==
1
)
)
)
begin
RXRDY
<=
!
CUARTOl0
;
end
end
end
end
end
endgenerate
always
@
(
posedge
CLK
or
negedge
CUARTI1
)
begin
if
(
(
!
CUARTI1
)
||
(
!
CUARTl1
)
)
begin
CUARTOO0
<=
1
'b
0
;
CUARTl1l
<=
1
'b
0
;
end
else
begin
CUARTl1l
<=
CUARTI1l
;
CUARTOO0
<=
CUARTl1l
;
end
end
always
@
(
posedge
CLK
or
negedge
CUARTI1
)
begin
if
(
(
!
CUARTI1
)
||
(
!
CUARTl1
)
)
begin
CUARTOI0
<=
1
'b
0
;
CUARTlO0
<=
1
'b
0
;
end
else
begin
CUARTlO0
<=
CUARTIO0
;
CUARTOI0
<=
CUARTlO0
;
end
end
always
@
(
posedge
CLK
or
negedge
CUARTI1
)
begin
if
(
(
!
CUARTI1
)
||
(
!
CUARTl1
)
)
begin
CUARTll0
<=
`CUARTOII
;
end
else
begin
CUARTll0
<=
CUARTO00
;
end
end
always
@
(
CUARTll0
,
CUARTOl0
,
CUARTlIl
)
begin
CUARTO00
=
CUARTll0
;
CUARTOll
=
1
'b
1
;
CUARTII0
=
1
'b
0
;
case
(
CUARTll0
)
`CUARTOII
:
if
(
CUARTOl0
==
1
'b
1
&&
CUARTlIl
==
1
'b
0
)
begin
CUARTO00
=
`CUARTIII
;
CUARTOll
=
1
'b
0
;
end
`CUARTIII
:
CUARTO00
=
`CUARTlII
;
`CUARTlII
:
CUARTO00
=
`CUARTOlI
;
`CUARTOlI
:
begin
CUARTO00
=
`CUARTOII
;
CUARTII0
=
1
'b
1
;
end
endcase
end
always
@
(
posedge
CLK
or
negedge
CUARTI1
)
begin
if
(
(
!
CUARTI1
)
||
(
!
CUARTl1
)
)
begin
CUARTIOl
<=
{
8
{
1
'b
0
}
}
;
end
else
begin
if
(
CUARTII0
==
1
'b
1
)
begin
CUARTIOl
<=
CUARTl1I
;
end
end
end
always
@
(
posedge
CLK
or
negedge
CUARTI1
)
begin
if
(
(
!
CUARTI1
)
||
(
!
CUARTl1
)
)
begin
CUARTOl0
<=
1
'b
1
;
CUARTIl0
<=
1
'b
1
;
end
else
begin
if
(
CUARTII0
==
1
'b
1
)
begin
CUARTOl0
<=
1
'b
0
;
end
else
begin
if
(
CSN
==
1
'b
0
&&
OEN
==
1
'b
0
)
begin
if
(
RX_FIFO
==
1
)
begin
if
(
!
PARITY_ERR
)
begin
CUARTOl0
<=
1
'b
1
;
end
end
else
begin
CUARTOl0
<=
1
'b
1
;
end
end
end
CUARTIl0
<=
CUARTOl0
;
end
end
always
@
(
posedge
CLK
or
negedge
CUARTI1
)
begin
if
(
(
!
CUARTI1
)
||
(
!
CUARTl1
)
)
begin
CUARTO10
<=
1
'b
0
;
end
else
begin
if
(
CUARTI0I
==
1
'b
0
&&
CUARTI0l
==
1
'b
1
)
CUARTO10
<=
1
'b
1
;
else
if
(
CUARTI10
==
1
'b
1
)
CUARTO10
<=
1
'b
0
;
else
CUARTO10
<=
CUARTO10
;
end
end
assign
OVERFLOW
=
(
RX_FIFO
==
1
'b
0
)
?
CUARTIlI
:
CUARTO10
;
assign
CUARTO0I
=
(
(
PARITY_ERR
==
1
'b
1
)
||
CUARTI0l
==
1
'b
1
)
?
1
'b
1
:
CUARTI0I
;
COREUART_C0_COREUART_C0_0_Clock_gen
#
(
.BAUD_VAL_FRCTN_EN
(
BAUD_VAL_FRCTN_EN
)
,
.SYNC_RESET
(
SYNC_RESET
)
)
CUARTOO1
(
.CUARTII
(
CLK
)
,
.CUARTlI
(
RESET_N
)
,
.CUARTOl
(
BAUD_VAL
)
,
.CUARTIl
(
CUARTIl
)
,
.CUARTll
(
CUARTll
)
,
.BAUD_VAL_FRACTION
(
BAUD_VAL_FRACTION
)
)
;
COREUART_C0_COREUART_C0_0_Tx_async
#
(
.TX_FIFO
(
TX_FIFO
)
,
.SYNC_RESET
(
SYNC_RESET
)
)
CUARTIO1
(
.CUARTII
(
CLK
)
,
.CUARTll
(
CUARTll
)
,
.CUARTlI
(
RESET_N
)
,
.CUARTl0I
(
CUARTl0I
)
,
.CUARTO1I
(
CUARTO1I
)
,
.CUARTI1I
(
CUARTI1I
)
,
.CUARTlO1
(
CUARTIIl
)
,
.CUARTOI1
(
CUARTO0l
)
,
.CUARTII1
(
BIT8
)
,
.CUARTlI1
(
PARITY_EN
)
,
.CUARTOl1
(
ODD_N_EVEN
)
,
.CUARTIl1
(
TXRDY
)
,
.CUARTll1
(
TX
)
,
.CUARTlll
(
CUARTlll
)
)
;
COREUART_C0_COREUART_C0_0_Rx_async
#
(
.RX_FIFO
(
RX_FIFO
)
,
.SYNC_RESET
(
SYNC_RESET
)
)
CUARTO01
(
.CUARTII
(
CLK
)
,
.CUARTIl
(
CUARTIl
)
,
.CUARTlI
(
RESET_N
)
,
.CUARTII1
(
BIT8
)
,
.CUARTlI1
(
PARITY_EN
)
,
.CUARTOl1
(
ODD_N_EVEN
)
,
.CUARTOOl
(
CUARTOOl
)
,
.CUARTl0l
(
CUARTl0l
)
,
.CUARTI01
(
FRAMING_ERR
)
,
.CUARTO1l
(
CUARTO1l
)
,
.CUARTI00
(
CUARTI00
)
,
.CUARTl00
(
CUARTl00
)
,
.CUARTl01
(
RX
)
,
.CUARTO11
(
CUARTIlI
)
,
.CUARTI11
(
PARITY_ERR
)
,
.CUARTI1l
(
CUARTI1l
)
,
.CUARTIO0
(
CUARTIO0
)
,
.CUARTllI
(
CUARTllI
)
,
.CUARTlOl
(
CUARTlOl
)
,
.CUARTI0I
(
CUARTI0I
)
)
;
generate
if
(
TX_FIFO
==
1
'b
1
)
begin
COREUART_C0_COREUART_C0_0_fifo_256x8
#
(
.SYNC_RESET
(
SYNC_RESET
)
)
CUARTl11
(
.CUARTOOOI
(
CUARTI1I
)
,
.CUARTIOOI
(
CLK
)
,
.CUARTlOOI
(
CLK
)
,
.CUARTOIOI
(
CUARTO1I
)
,
.WRB
(
CUARTIll
)
,
.RDB
(
CUARTlll
)
,
.RESET
(
RESET_N
)
,
.FULL
(
CUARTO0l
)
,
.EMPTY
(
CUARTIIl
)
)
;
end
else
begin
assign
CUARTO0l
=
1
'b
0
;
assign
CUARTIIl
=
1
'b
0
;
assign
CUARTI1I
=
8
'b
0
;
end
endgenerate
generate
if
(
RX_FIFO
==
1
'b
1
)
begin
COREUART_C0_COREUART_C0_0_fifo_256x8
#
(
.SYNC_RESET
(
SYNC_RESET
)
)
CUARTIIOI
(
.CUARTOOOI
(
CUARTl1I
)
,
.CUARTIOOI
(
CLK
)
,
.CUARTlOOI
(
CLK
)
,
.CUARTOIOI
(
CUARTOIl
)
,
.WRB
(
CUARTO0I
)
,
.RDB
(
CUARTOll
)
,
.RESET
(
RESET_N
)
,
.FULL
(
CUARTI0l
)
,
.EMPTY
(
CUARTlIl
)
)
;
end
else
begin
assign
CUARTI0l
=
1
'b
0
;
assign
CUARTlIl
=
1
'b
0
;
assign
CUARTl1I
=
8
'b
0
;
end
endgenerate
endmodule
